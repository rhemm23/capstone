module ctrl_test;


endmodule
