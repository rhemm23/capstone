module ctrl_test;


reg clk, rst_n;


ctrl_unit ctrlUnit(.*);

endmodule
