module iru_cos_lut
  (
    /*
     * Inputs
     */
    input [5:0] d,

    /*
     * Outputs
     */
    output reg [8:0] q
  );

  always_comb begin
    case (d)
      9'b000000: q <= 8'b010000000;
      9'b000001: q <= 8'b001111110;
      9'b000010: q <= 8'b001111000;
      9'b000011: q <= 8'b001101110;
      9'b000100: q <= 8'b001100010;
      9'b000101: q <= 8'b001010010;
      9'b000110: q <= 8'b001000000;
      9'b000111: q <= 8'b000101011;
      9'b001000: q <= 8'b000010110;
      9'b001001: q <= 8'b000000000;
      9'b001010: q <= 8'b100010110;
      9'b001011: q <= 8'b100101011;
      9'b001100: q <= 8'b100111111;
      9'b001101: q <= 8'b101010010;
      9'b001110: q <= 8'b101100010;
      9'b001111: q <= 8'b101101110;
      9'b010000: q <= 8'b101111000;
      9'b010001: q <= 8'b101111110;
      9'b010010: q <= 8'b110000000;
      9'b010011: q <= 8'b101111110;
      9'b010100: q <= 8'b101111000;
      9'b010101: q <= 8'b101101110;
      9'b010110: q <= 8'b101100010;
      9'b010111: q <= 8'b101010010;
      9'b011000: q <= 8'b101000000;
      9'b011001: q <= 8'b100101011;
      9'b011010: q <= 8'b100010110;
      9'b011011: q <= 8'b100000000;
      9'b011100: q <= 8'b000010110;
      9'b011101: q <= 8'b000101011;
      9'b011110: q <= 8'b001000000;
      9'b011111: q <= 8'b001010010;
      9'b100000: q <= 8'b001100010;
      9'b100001: q <= 8'b001101110;
      9'b100010: q <= 8'b001111000;
      9'b100011: q <= 8'b001111110;
      default: q <= 0;
    endcase
  end

endmodule
