module pipeline_wrapper
(

);

endmodule