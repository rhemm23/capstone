`ifndef MEM_TYPES_VH
`define MEM_TYPES_VH

import mem_types::*;

`endif
