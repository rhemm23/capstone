`ifndef DATA_TYPES_VH
`define DATA_TYPES_VH

import data_types::*;

`endif
