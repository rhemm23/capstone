module ipgu_mult_lut
  (
    /*
     * Inputs
     */
    input [2:0] scaleNum,//which downscale ratio to use/multiplier
    input [8:0] addr,//9 bits for addr

    /*
     * Outputs
     */
    output wire [8:0] addrOut
  );

  reg [8:0] q [5];
  always_comb begin
    case (addr[9-1:0])
      9'b000000000: q[0] <= 9'b000000000;
      9'b000000001: q[0] <= 9'b000000000;
      9'b000000010: q[0] <= 9'b000000001;
      9'b000000011: q[0] <= 9'b000000010;
      9'b000000100: q[0] <= 9'b000000011;
      9'b000000101: q[0] <= 9'b000000100;
      9'b000000110: q[0] <= 9'b000000100;
      9'b000000111: q[0] <= 9'b000000101;
      9'b000001000: q[0] <= 9'b000000110;
      9'b000001001: q[0] <= 9'b000000111;
      9'b000001010: q[0] <= 9'b000001000;
      9'b000001011: q[0] <= 9'b000001000;
      9'b000001100: q[0] <= 9'b000001001;
      9'b000001101: q[0] <= 9'b000001010;
      9'b000001110: q[0] <= 9'b000001011;
      9'b000001111: q[0] <= 9'b000001100;
      9'b000010000: q[0] <= 9'b000001100;
      9'b000010001: q[0] <= 9'b000001101;
      9'b000010010: q[0] <= 9'b000001110;
      9'b000010011: q[0] <= 9'b000001111;
      9'b000010100: q[0] <= 9'b000010000;
      9'b000010101: q[0] <= 9'b000010000;
      9'b000010110: q[0] <= 9'b000010001;
      9'b000010111: q[0] <= 9'b000010010;
      9'b000011000: q[0] <= 9'b000010011;
      9'b000011001: q[0] <= 9'b000010100;
      9'b000011010: q[0] <= 9'b000010100;
      9'b000011011: q[0] <= 9'b000010101;
      9'b000011100: q[0] <= 9'b000010110;
      9'b000011101: q[0] <= 9'b000010111;
      9'b000011110: q[0] <= 9'b000011000;
      9'b000011111: q[0] <= 9'b000011000;
      9'b000100000: q[0] <= 9'b000011001;
      9'b000100001: q[0] <= 9'b000011010;
      9'b000100010: q[0] <= 9'b000011011;
      9'b000100011: q[0] <= 9'b000011100;
      9'b000100100: q[0] <= 9'b000011100;
      9'b000100101: q[0] <= 9'b000011101;
      9'b000100110: q[0] <= 9'b000011110;
      9'b000100111: q[0] <= 9'b000011111;
      9'b000101000: q[0] <= 9'b000100000;
      9'b000101001: q[0] <= 9'b000100000;
      9'b000101010: q[0] <= 9'b000100001;
      9'b000101011: q[0] <= 9'b000100010;
      9'b000101100: q[0] <= 9'b000100011;
      9'b000101101: q[0] <= 9'b000100100;
      9'b000101110: q[0] <= 9'b000100100;
      9'b000101111: q[0] <= 9'b000100101;
      9'b000110000: q[0] <= 9'b000100110;
      9'b000110001: q[0] <= 9'b000100111;
      9'b000110010: q[0] <= 9'b000101000;
      9'b000110011: q[0] <= 9'b000101000;
      9'b000110100: q[0] <= 9'b000101001;
      9'b000110101: q[0] <= 9'b000101010;
      9'b000110110: q[0] <= 9'b000101011;
      9'b000110111: q[0] <= 9'b000101100;
      9'b000111000: q[0] <= 9'b000101100;
      9'b000111001: q[0] <= 9'b000101101;
      9'b000111010: q[0] <= 9'b000101110;
      9'b000111011: q[0] <= 9'b000101111;
      9'b000111100: q[0] <= 9'b000110000;
      9'b000111101: q[0] <= 9'b000110000;
      9'b000111110: q[0] <= 9'b000110001;
      9'b000111111: q[0] <= 9'b000110010;
      9'b001000000: q[0] <= 9'b000110011;
      9'b001000001: q[0] <= 9'b000110100;
      9'b001000010: q[0] <= 9'b000110100;
      9'b001000011: q[0] <= 9'b000110101;
      9'b001000100: q[0] <= 9'b000110110;
      9'b001000101: q[0] <= 9'b000110111;
      9'b001000110: q[0] <= 9'b000111000;
      9'b001000111: q[0] <= 9'b000111000;
      9'b001001000: q[0] <= 9'b000111001;
      9'b001001001: q[0] <= 9'b000111010;
      9'b001001010: q[0] <= 9'b000111011;
      9'b001001011: q[0] <= 9'b000111100;
      9'b001001100: q[0] <= 9'b000111100;
      9'b001001101: q[0] <= 9'b000111101;
      9'b001001110: q[0] <= 9'b000111110;
      9'b001001111: q[0] <= 9'b000111111;
      9'b001010000: q[0] <= 9'b001000000;
      9'b001010001: q[0] <= 9'b001000000;
      9'b001010010: q[0] <= 9'b001000001;
      9'b001010011: q[0] <= 9'b001000010;
      9'b001010100: q[0] <= 9'b001000011;
      9'b001010101: q[0] <= 9'b001000100;
      9'b001010110: q[0] <= 9'b001000100;
      9'b001010111: q[0] <= 9'b001000101;
      9'b001011000: q[0] <= 9'b001000110;
      9'b001011001: q[0] <= 9'b001000111;
      9'b001011010: q[0] <= 9'b001001000;
      9'b001011011: q[0] <= 9'b001001000;
      9'b001011100: q[0] <= 9'b001001001;
      9'b001011101: q[0] <= 9'b001001010;
      9'b001011110: q[0] <= 9'b001001011;
      9'b001011111: q[0] <= 9'b001001100;
      9'b001100000: q[0] <= 9'b001001100;
      9'b001100001: q[0] <= 9'b001001101;
      9'b001100010: q[0] <= 9'b001001110;
      9'b001100011: q[0] <= 9'b001001111;
      9'b001100100: q[0] <= 9'b001010000;
      9'b001100101: q[0] <= 9'b001010000;
      9'b001100110: q[0] <= 9'b001010001;
      9'b001100111: q[0] <= 9'b001010010;
      9'b001101000: q[0] <= 9'b001010011;
      9'b001101001: q[0] <= 9'b001010100;
      9'b001101010: q[0] <= 9'b001010100;
      9'b001101011: q[0] <= 9'b001010101;
      9'b001101100: q[0] <= 9'b001010110;
      9'b001101101: q[0] <= 9'b001010111;
      9'b001101110: q[0] <= 9'b001011000;
      9'b001101111: q[0] <= 9'b001011000;
      9'b001110000: q[0] <= 9'b001011001;
      9'b001110001: q[0] <= 9'b001011010;
      9'b001110010: q[0] <= 9'b001011011;
      9'b001110011: q[0] <= 9'b001011100;
      9'b001110100: q[0] <= 9'b001011100;
      9'b001110101: q[0] <= 9'b001011101;
      9'b001110110: q[0] <= 9'b001011110;
      9'b001110111: q[0] <= 9'b001011111;
      9'b001111000: q[0] <= 9'b001100000;
      9'b001111001: q[0] <= 9'b001100000;
      9'b001111010: q[0] <= 9'b001100001;
      9'b001111011: q[0] <= 9'b001100010;
      9'b001111100: q[0] <= 9'b001100011;
      9'b001111101: q[0] <= 9'b001100100;
      9'b001111110: q[0] <= 9'b001100100;
      9'b001111111: q[0] <= 9'b001100101;
      9'b010000000: q[0] <= 9'b001100110;
      9'b010000001: q[0] <= 9'b001100111;
      9'b010000010: q[0] <= 9'b001101000;
      9'b010000011: q[0] <= 9'b001101000;
      9'b010000100: q[0] <= 9'b001101001;
      9'b010000101: q[0] <= 9'b001101010;
      9'b010000110: q[0] <= 9'b001101011;
      9'b010000111: q[0] <= 9'b001101100;
      9'b010001000: q[0] <= 9'b001101100;
      9'b010001001: q[0] <= 9'b001101101;
      9'b010001010: q[0] <= 9'b001101110;
      9'b010001011: q[0] <= 9'b001101111;
      9'b010001100: q[0] <= 9'b001110000;
      9'b010001101: q[0] <= 9'b001110000;
      9'b010001110: q[0] <= 9'b001110001;
      9'b010001111: q[0] <= 9'b001110010;
      9'b010010000: q[0] <= 9'b001110011;
      9'b010010001: q[0] <= 9'b001110100;
      9'b010010010: q[0] <= 9'b001110100;
      9'b010010011: q[0] <= 9'b001110101;
      9'b010010100: q[0] <= 9'b001110110;
      9'b010010101: q[0] <= 9'b001110111;
      9'b010010110: q[0] <= 9'b001111000;
      9'b010010111: q[0] <= 9'b001111000;
      9'b010011000: q[0] <= 9'b001111001;
      9'b010011001: q[0] <= 9'b001111010;
      9'b010011010: q[0] <= 9'b001111011;
      9'b010011011: q[0] <= 9'b001111100;
      9'b010011100: q[0] <= 9'b001111100;
      9'b010011101: q[0] <= 9'b001111101;
      9'b010011110: q[0] <= 9'b001111110;
      9'b010011111: q[0] <= 9'b001111111;
      9'b010100000: q[0] <= 9'b010000000;
      9'b010100001: q[0] <= 9'b010000000;
      9'b010100010: q[0] <= 9'b010000001;
      9'b010100011: q[0] <= 9'b010000010;
      9'b010100100: q[0] <= 9'b010000011;
      9'b010100101: q[0] <= 9'b010000100;
      9'b010100110: q[0] <= 9'b010000100;
      9'b010100111: q[0] <= 9'b010000101;
      9'b010101000: q[0] <= 9'b010000110;
      9'b010101001: q[0] <= 9'b010000111;
      9'b010101010: q[0] <= 9'b010001000;
      9'b010101011: q[0] <= 9'b010001000;
      9'b010101100: q[0] <= 9'b010001001;
      9'b010101101: q[0] <= 9'b010001010;
      9'b010101110: q[0] <= 9'b010001011;
      9'b010101111: q[0] <= 9'b010001100;
      9'b010110000: q[0] <= 9'b010001100;
      9'b010110001: q[0] <= 9'b010001101;
      9'b010110010: q[0] <= 9'b010001110;
      9'b010110011: q[0] <= 9'b010001111;
      9'b010110100: q[0] <= 9'b010010000;
      9'b010110101: q[0] <= 9'b010010000;
      9'b010110110: q[0] <= 9'b010010001;
      9'b010110111: q[0] <= 9'b010010010;
      9'b010111000: q[0] <= 9'b010010011;
      9'b010111001: q[0] <= 9'b010010100;
      9'b010111010: q[0] <= 9'b010010100;
      9'b010111011: q[0] <= 9'b010010101;
      9'b010111100: q[0] <= 9'b010010110;
      9'b010111101: q[0] <= 9'b010010111;
      9'b010111110: q[0] <= 9'b010011000;
      9'b010111111: q[0] <= 9'b010011000;
      9'b011000000: q[0] <= 9'b010011001;
      9'b011000001: q[0] <= 9'b010011010;
      9'b011000010: q[0] <= 9'b010011011;
      9'b011000011: q[0] <= 9'b010011100;
      9'b011000100: q[0] <= 9'b010011100;
      9'b011000101: q[0] <= 9'b010011101;
      9'b011000110: q[0] <= 9'b010011110;
      9'b011000111: q[0] <= 9'b010011111;
      9'b011001000: q[0] <= 9'b010100000;
      9'b011001001: q[0] <= 9'b010100000;
      9'b011001010: q[0] <= 9'b010100001;
      9'b011001011: q[0] <= 9'b010100010;
      9'b011001100: q[0] <= 9'b010100011;
      9'b011001101: q[0] <= 9'b010100100;
      9'b011001110: q[0] <= 9'b010100100;
      9'b011001111: q[0] <= 9'b010100101;
      9'b011010000: q[0] <= 9'b010100110;
      9'b011010001: q[0] <= 9'b010100111;
      9'b011010010: q[0] <= 9'b010101000;
      9'b011010011: q[0] <= 9'b010101000;
      9'b011010100: q[0] <= 9'b010101001;
      9'b011010101: q[0] <= 9'b010101010;
      9'b011010110: q[0] <= 9'b010101011;
      9'b011010111: q[0] <= 9'b010101100;
      9'b011011000: q[0] <= 9'b010101100;
      9'b011011001: q[0] <= 9'b010101101;
      9'b011011010: q[0] <= 9'b010101110;
      9'b011011011: q[0] <= 9'b010101111;
      9'b011011100: q[0] <= 9'b010110000;
      9'b011011101: q[0] <= 9'b010110000;
      9'b011011110: q[0] <= 9'b010110001;
      9'b011011111: q[0] <= 9'b010110010;
      9'b011100000: q[0] <= 9'b010110011;
      9'b011100001: q[0] <= 9'b010110100;
      9'b011100010: q[0] <= 9'b010110100;
      9'b011100011: q[0] <= 9'b010110101;
      9'b011100100: q[0] <= 9'b010110110;
      9'b011100101: q[0] <= 9'b010110111;
      9'b011100110: q[0] <= 9'b010111000;
      9'b011100111: q[0] <= 9'b010111000;
      9'b011101000: q[0] <= 9'b010111001;
      9'b011101001: q[0] <= 9'b010111010;
      9'b011101010: q[0] <= 9'b010111011;
      9'b011101011: q[0] <= 9'b010111100;
      9'b011101100: q[0] <= 9'b010111100;
      9'b011101101: q[0] <= 9'b010111101;
      9'b011101110: q[0] <= 9'b010111110;
      9'b011101111: q[0] <= 9'b010111111;
      9'b011110000: q[0] <= 9'b011000000;
      9'b011110001: q[0] <= 9'b011000000;
      9'b011110010: q[0] <= 9'b011000001;
      9'b011110011: q[0] <= 9'b011000010;
      9'b011110100: q[0] <= 9'b011000011;
      9'b011110101: q[0] <= 9'b011000100;
      9'b011110110: q[0] <= 9'b011000100;
      9'b011110111: q[0] <= 9'b011000101;
      9'b011111000: q[0] <= 9'b011000110;
      9'b011111001: q[0] <= 9'b011000111;
      9'b011111010: q[0] <= 9'b011001000;
      9'b011111011: q[0] <= 9'b011001000;
      9'b011111100: q[0] <= 9'b011001001;
      9'b011111101: q[0] <= 9'b011001010;
      9'b011111110: q[0] <= 9'b011001011;
      9'b011111111: q[0] <= 9'b011001100;
      9'b100000000: q[0] <= 9'b011001100;
      9'b100000001: q[0] <= 9'b011001101;
      9'b100000010: q[0] <= 9'b011001110;
      9'b100000011: q[0] <= 9'b011001111;
      9'b100000100: q[0] <= 9'b011010000;
      9'b100000101: q[0] <= 9'b011010000;
      9'b100000110: q[0] <= 9'b011010001;
      9'b100000111: q[0] <= 9'b011010010;
      9'b100001000: q[0] <= 9'b011010011;
      9'b100001001: q[0] <= 9'b011010100;
      9'b100001010: q[0] <= 9'b011010100;
      9'b100001011: q[0] <= 9'b011010101;
      9'b100001100: q[0] <= 9'b011010110;
      9'b100001101: q[0] <= 9'b011010111;
      9'b100001110: q[0] <= 9'b011011000;
      9'b100001111: q[0] <= 9'b011011000;
      9'b100010000: q[0] <= 9'b011011001;
      9'b100010001: q[0] <= 9'b011011010;
      9'b100010010: q[0] <= 9'b011011011;
      9'b100010011: q[0] <= 9'b011011100;
      9'b100010100: q[0] <= 9'b011011100;
      9'b100010101: q[0] <= 9'b011011101;
      9'b100010110: q[0] <= 9'b011011110;
      9'b100010111: q[0] <= 9'b011011111;
      9'b100011000: q[0] <= 9'b011100000;
      9'b100011001: q[0] <= 9'b011100000;
      9'b100011010: q[0] <= 9'b011100001;
      9'b100011011: q[0] <= 9'b011100010;
      9'b100011100: q[0] <= 9'b011100011;
      9'b100011101: q[0] <= 9'b011100100;
      9'b100011110: q[0] <= 9'b011100100;
      9'b100011111: q[0] <= 9'b011100101;
      9'b100100000: q[0] <= 9'b011100110;
      9'b100100001: q[0] <= 9'b011100111;
      9'b100100010: q[0] <= 9'b011101000;
      9'b100100011: q[0] <= 9'b011101000;
      9'b100100100: q[0] <= 9'b011101001;
      9'b100100101: q[0] <= 9'b011101010;
      9'b100100110: q[0] <= 9'b011101011;
      9'b100100111: q[0] <= 9'b011101100;
      9'b100101000: q[0] <= 9'b011101100;
      9'b100101001: q[0] <= 9'b011101101;
      9'b100101010: q[0] <= 9'b011101110;
      9'b100101011: q[0] <= 9'b011101111;
      default: q[0] <= '0;
    endcase
    case (addr[8-1:0])
      8'b00000000: q[1] <= 9'b000000000;
      8'b00000001: q[1] <= 9'b000000000;
      8'b00000010: q[1] <= 9'b000000001;
      8'b00000011: q[1] <= 9'b000000010;
      8'b00000100: q[1] <= 9'b000000011;
      8'b00000101: q[1] <= 9'b000000011;
      8'b00000110: q[1] <= 9'b000000100;
      8'b00000111: q[1] <= 9'b000000101;
      8'b00001000: q[1] <= 9'b000000110;
      8'b00001001: q[1] <= 9'b000000110;
      8'b00001010: q[1] <= 9'b000000111;
      8'b00001011: q[1] <= 9'b000001000;
      8'b00001100: q[1] <= 9'b000001001;
      8'b00001101: q[1] <= 9'b000001001;
      8'b00001110: q[1] <= 9'b000001010;
      8'b00001111: q[1] <= 9'b000001011;
      8'b00010000: q[1] <= 9'b000001100;
      8'b00010001: q[1] <= 9'b000001100;
      8'b00010010: q[1] <= 9'b000001101;
      8'b00010011: q[1] <= 9'b000001110;
      8'b00010100: q[1] <= 9'b000001111;
      8'b00010101: q[1] <= 9'b000001111;
      8'b00010110: q[1] <= 9'b000010000;
      8'b00010111: q[1] <= 9'b000010001;
      8'b00011000: q[1] <= 9'b000010010;
      8'b00011001: q[1] <= 9'b000010010;
      8'b00011010: q[1] <= 9'b000010011;
      8'b00011011: q[1] <= 9'b000010100;
      8'b00011100: q[1] <= 9'b000010101;
      8'b00011101: q[1] <= 9'b000010101;
      8'b00011110: q[1] <= 9'b000010110;
      8'b00011111: q[1] <= 9'b000010111;
      8'b00100000: q[1] <= 9'b000011000;
      8'b00100001: q[1] <= 9'b000011000;
      8'b00100010: q[1] <= 9'b000011001;
      8'b00100011: q[1] <= 9'b000011010;
      8'b00100100: q[1] <= 9'b000011011;
      8'b00100101: q[1] <= 9'b000011011;
      8'b00100110: q[1] <= 9'b000011100;
      8'b00100111: q[1] <= 9'b000011101;
      8'b00101000: q[1] <= 9'b000011110;
      8'b00101001: q[1] <= 9'b000011110;
      8'b00101010: q[1] <= 9'b000011111;
      8'b00101011: q[1] <= 9'b000100000;
      8'b00101100: q[1] <= 9'b000100001;
      8'b00101101: q[1] <= 9'b000100001;
      8'b00101110: q[1] <= 9'b000100010;
      8'b00101111: q[1] <= 9'b000100011;
      8'b00110000: q[1] <= 9'b000100100;
      8'b00110001: q[1] <= 9'b000100100;
      8'b00110010: q[1] <= 9'b000100101;
      8'b00110011: q[1] <= 9'b000100110;
      8'b00110100: q[1] <= 9'b000100111;
      8'b00110101: q[1] <= 9'b000100111;
      8'b00110110: q[1] <= 9'b000101000;
      8'b00110111: q[1] <= 9'b000101001;
      8'b00111000: q[1] <= 9'b000101010;
      8'b00111001: q[1] <= 9'b000101010;
      8'b00111010: q[1] <= 9'b000101011;
      8'b00111011: q[1] <= 9'b000101100;
      8'b00111100: q[1] <= 9'b000101101;
      8'b00111101: q[1] <= 9'b000101101;
      8'b00111110: q[1] <= 9'b000101110;
      8'b00111111: q[1] <= 9'b000101111;
      8'b01000000: q[1] <= 9'b000110000;
      8'b01000001: q[1] <= 9'b000110000;
      8'b01000010: q[1] <= 9'b000110001;
      8'b01000011: q[1] <= 9'b000110010;
      8'b01000100: q[1] <= 9'b000110011;
      8'b01000101: q[1] <= 9'b000110011;
      8'b01000110: q[1] <= 9'b000110100;
      8'b01000111: q[1] <= 9'b000110101;
      8'b01001000: q[1] <= 9'b000110110;
      8'b01001001: q[1] <= 9'b000110110;
      8'b01001010: q[1] <= 9'b000110111;
      8'b01001011: q[1] <= 9'b000111000;
      8'b01001100: q[1] <= 9'b000111001;
      8'b01001101: q[1] <= 9'b000111001;
      8'b01001110: q[1] <= 9'b000111010;
      8'b01001111: q[1] <= 9'b000111011;
      8'b01010000: q[1] <= 9'b000111100;
      8'b01010001: q[1] <= 9'b000111100;
      8'b01010010: q[1] <= 9'b000111101;
      8'b01010011: q[1] <= 9'b000111110;
      8'b01010100: q[1] <= 9'b000111111;
      8'b01010101: q[1] <= 9'b000111111;
      8'b01010110: q[1] <= 9'b001000000;
      8'b01010111: q[1] <= 9'b001000001;
      8'b01011000: q[1] <= 9'b001000010;
      8'b01011001: q[1] <= 9'b001000010;
      8'b01011010: q[1] <= 9'b001000011;
      8'b01011011: q[1] <= 9'b001000100;
      8'b01011100: q[1] <= 9'b001000101;
      8'b01011101: q[1] <= 9'b001000101;
      8'b01011110: q[1] <= 9'b001000110;
      8'b01011111: q[1] <= 9'b001000111;
      8'b01100000: q[1] <= 9'b001001000;
      8'b01100001: q[1] <= 9'b001001000;
      8'b01100010: q[1] <= 9'b001001001;
      8'b01100011: q[1] <= 9'b001001010;
      8'b01100100: q[1] <= 9'b001001011;
      8'b01100101: q[1] <= 9'b001001011;
      8'b01100110: q[1] <= 9'b001001100;
      8'b01100111: q[1] <= 9'b001001101;
      8'b01101000: q[1] <= 9'b001001110;
      8'b01101001: q[1] <= 9'b001001110;
      8'b01101010: q[1] <= 9'b001001111;
      8'b01101011: q[1] <= 9'b001010000;
      8'b01101100: q[1] <= 9'b001010001;
      8'b01101101: q[1] <= 9'b001010001;
      8'b01101110: q[1] <= 9'b001010010;
      8'b01101111: q[1] <= 9'b001010011;
      8'b01110000: q[1] <= 9'b001010100;
      8'b01110001: q[1] <= 9'b001010100;
      8'b01110010: q[1] <= 9'b001010101;
      8'b01110011: q[1] <= 9'b001010110;
      8'b01110100: q[1] <= 9'b001010111;
      8'b01110101: q[1] <= 9'b001010111;
      8'b01110110: q[1] <= 9'b001011000;
      8'b01110111: q[1] <= 9'b001011001;
      8'b01111000: q[1] <= 9'b001011010;
      8'b01111001: q[1] <= 9'b001011010;
      8'b01111010: q[1] <= 9'b001011011;
      8'b01111011: q[1] <= 9'b001011100;
      8'b01111100: q[1] <= 9'b001011101;
      8'b01111101: q[1] <= 9'b001011101;
      8'b01111110: q[1] <= 9'b001011110;
      8'b01111111: q[1] <= 9'b001011111;
      8'b10000000: q[1] <= 9'b001100000;
      8'b10000001: q[1] <= 9'b001100000;
      8'b10000010: q[1] <= 9'b001100001;
      8'b10000011: q[1] <= 9'b001100010;
      8'b10000100: q[1] <= 9'b001100011;
      8'b10000101: q[1] <= 9'b001100011;
      8'b10000110: q[1] <= 9'b001100100;
      8'b10000111: q[1] <= 9'b001100101;
      8'b10001000: q[1] <= 9'b001100110;
      8'b10001001: q[1] <= 9'b001100110;
      8'b10001010: q[1] <= 9'b001100111;
      8'b10001011: q[1] <= 9'b001101000;
      8'b10001100: q[1] <= 9'b001101001;
      8'b10001101: q[1] <= 9'b001101001;
      8'b10001110: q[1] <= 9'b001101010;
      8'b10001111: q[1] <= 9'b001101011;
      8'b10010000: q[1] <= 9'b001101100;
      8'b10010001: q[1] <= 9'b001101100;
      8'b10010010: q[1] <= 9'b001101101;
      8'b10010011: q[1] <= 9'b001101110;
      8'b10010100: q[1] <= 9'b001101111;
      8'b10010101: q[1] <= 9'b001101111;
      8'b10010110: q[1] <= 9'b001110000;
      8'b10010111: q[1] <= 9'b001110001;
      8'b10011000: q[1] <= 9'b001110010;
      8'b10011001: q[1] <= 9'b001110010;
      8'b10011010: q[1] <= 9'b001110011;
      8'b10011011: q[1] <= 9'b001110100;
      8'b10011100: q[1] <= 9'b001110101;
      8'b10011101: q[1] <= 9'b001110101;
      8'b10011110: q[1] <= 9'b001110110;
      8'b10011111: q[1] <= 9'b001110111;
      8'b10100000: q[1] <= 9'b001111000;
      8'b10100001: q[1] <= 9'b001111000;
      8'b10100010: q[1] <= 9'b001111001;
      8'b10100011: q[1] <= 9'b001111010;
      8'b10100100: q[1] <= 9'b001111011;
      8'b10100101: q[1] <= 9'b001111011;
      8'b10100110: q[1] <= 9'b001111100;
      8'b10100111: q[1] <= 9'b001111101;
      8'b10101000: q[1] <= 9'b001111110;
      8'b10101001: q[1] <= 9'b001111110;
      8'b10101010: q[1] <= 9'b001111111;
      8'b10101011: q[1] <= 9'b010000000;
      8'b10101100: q[1] <= 9'b010000001;
      8'b10101101: q[1] <= 9'b010000001;
      8'b10101110: q[1] <= 9'b010000010;
      8'b10101111: q[1] <= 9'b010000011;
      8'b10110000: q[1] <= 9'b010000100;
      8'b10110001: q[1] <= 9'b010000100;
      8'b10110010: q[1] <= 9'b010000101;
      8'b10110011: q[1] <= 9'b010000110;
      8'b10110100: q[1] <= 9'b010000111;
      8'b10110101: q[1] <= 9'b010000111;
      8'b10110110: q[1] <= 9'b010001000;
      8'b10110111: q[1] <= 9'b010001001;
      8'b10111000: q[1] <= 9'b010001010;
      8'b10111001: q[1] <= 9'b010001010;
      8'b10111010: q[1] <= 9'b010001011;
      8'b10111011: q[1] <= 9'b010001100;
      8'b10111100: q[1] <= 9'b010001101;
      8'b10111101: q[1] <= 9'b010001101;
      8'b10111110: q[1] <= 9'b010001110;
      8'b10111111: q[1] <= 9'b010001111;
      8'b11000000: q[1] <= 9'b010010000;
      8'b11000001: q[1] <= 9'b010010000;
      8'b11000010: q[1] <= 9'b010010001;
      8'b11000011: q[1] <= 9'b010010010;
      8'b11000100: q[1] <= 9'b010010011;
      8'b11000101: q[1] <= 9'b010010011;
      8'b11000110: q[1] <= 9'b010010100;
      8'b11000111: q[1] <= 9'b010010101;
      8'b11001000: q[1] <= 9'b010010110;
      8'b11001001: q[1] <= 9'b010010110;
      8'b11001010: q[1] <= 9'b010010111;
      8'b11001011: q[1] <= 9'b010011000;
      8'b11001100: q[1] <= 9'b010011001;
      8'b11001101: q[1] <= 9'b010011001;
      8'b11001110: q[1] <= 9'b010011010;
      8'b11001111: q[1] <= 9'b010011011;
      8'b11010000: q[1] <= 9'b010011100;
      8'b11010001: q[1] <= 9'b010011100;
      8'b11010010: q[1] <= 9'b010011101;
      8'b11010011: q[1] <= 9'b010011110;
      8'b11010100: q[1] <= 9'b010011111;
      8'b11010101: q[1] <= 9'b010011111;
      8'b11010110: q[1] <= 9'b010100000;
      8'b11010111: q[1] <= 9'b010100001;
      8'b11011000: q[1] <= 9'b010100010;
      8'b11011001: q[1] <= 9'b010100010;
      8'b11011010: q[1] <= 9'b010100011;
      8'b11011011: q[1] <= 9'b010100100;
      8'b11011100: q[1] <= 9'b010100101;
      8'b11011101: q[1] <= 9'b010100101;
      8'b11011110: q[1] <= 9'b010100110;
      8'b11011111: q[1] <= 9'b010100111;
      8'b11100000: q[1] <= 9'b010101000;
      8'b11100001: q[1] <= 9'b010101000;
      8'b11100010: q[1] <= 9'b010101001;
      8'b11100011: q[1] <= 9'b010101010;
      8'b11100100: q[1] <= 9'b010101011;
      8'b11100101: q[1] <= 9'b010101011;
      8'b11100110: q[1] <= 9'b010101100;
      8'b11100111: q[1] <= 9'b010101101;
      8'b11101000: q[1] <= 9'b010101110;
      8'b11101001: q[1] <= 9'b010101110;
      8'b11101010: q[1] <= 9'b010101111;
      8'b11101011: q[1] <= 9'b010110000;
      8'b11101100: q[1] <= 9'b010110001;
      8'b11101101: q[1] <= 9'b010110001;
      8'b11101110: q[1] <= 9'b010110010;
      8'b11101111: q[1] <= 9'b010110011;
      default: q[1] <= '0;
    endcase
    case (addr[8-1:0])
      8'b00000000: q[2] <= 9'b000000000;
      8'b00000001: q[2] <= 9'b000000000;
      8'b00000010: q[2] <= 9'b000000001;
      8'b00000011: q[2] <= 9'b000000010;
      8'b00000100: q[2] <= 9'b000000010;
      8'b00000101: q[2] <= 9'b000000011;
      8'b00000110: q[2] <= 9'b000000100;
      8'b00000111: q[2] <= 9'b000000100;
      8'b00001000: q[2] <= 9'b000000101;
      8'b00001001: q[2] <= 9'b000000110;
      8'b00001010: q[2] <= 9'b000000110;
      8'b00001011: q[2] <= 9'b000000111;
      8'b00001100: q[2] <= 9'b000001000;
      8'b00001101: q[2] <= 9'b000001000;
      8'b00001110: q[2] <= 9'b000001001;
      8'b00001111: q[2] <= 9'b000001010;
      8'b00010000: q[2] <= 9'b000001010;
      8'b00010001: q[2] <= 9'b000001011;
      8'b00010010: q[2] <= 9'b000001100;
      8'b00010011: q[2] <= 9'b000001100;
      8'b00010100: q[2] <= 9'b000001101;
      8'b00010101: q[2] <= 9'b000001110;
      8'b00010110: q[2] <= 9'b000001110;
      8'b00010111: q[2] <= 9'b000001111;
      8'b00011000: q[2] <= 9'b000010000;
      8'b00011001: q[2] <= 9'b000010000;
      8'b00011010: q[2] <= 9'b000010001;
      8'b00011011: q[2] <= 9'b000010010;
      8'b00011100: q[2] <= 9'b000010010;
      8'b00011101: q[2] <= 9'b000010011;
      8'b00011110: q[2] <= 9'b000010100;
      8'b00011111: q[2] <= 9'b000010100;
      8'b00100000: q[2] <= 9'b000010101;
      8'b00100001: q[2] <= 9'b000010110;
      8'b00100010: q[2] <= 9'b000010110;
      8'b00100011: q[2] <= 9'b000010111;
      8'b00100100: q[2] <= 9'b000011000;
      8'b00100101: q[2] <= 9'b000011000;
      8'b00100110: q[2] <= 9'b000011001;
      8'b00100111: q[2] <= 9'b000011010;
      8'b00101000: q[2] <= 9'b000011010;
      8'b00101001: q[2] <= 9'b000011011;
      8'b00101010: q[2] <= 9'b000011100;
      8'b00101011: q[2] <= 9'b000011100;
      8'b00101100: q[2] <= 9'b000011101;
      8'b00101101: q[2] <= 9'b000011110;
      8'b00101110: q[2] <= 9'b000011110;
      8'b00101111: q[2] <= 9'b000011111;
      8'b00110000: q[2] <= 9'b000100000;
      8'b00110001: q[2] <= 9'b000100000;
      8'b00110010: q[2] <= 9'b000100001;
      8'b00110011: q[2] <= 9'b000100010;
      8'b00110100: q[2] <= 9'b000100010;
      8'b00110101: q[2] <= 9'b000100011;
      8'b00110110: q[2] <= 9'b000100100;
      8'b00110111: q[2] <= 9'b000100100;
      8'b00111000: q[2] <= 9'b000100101;
      8'b00111001: q[2] <= 9'b000100110;
      8'b00111010: q[2] <= 9'b000100110;
      8'b00111011: q[2] <= 9'b000100111;
      8'b00111100: q[2] <= 9'b000101000;
      8'b00111101: q[2] <= 9'b000101000;
      8'b00111110: q[2] <= 9'b000101001;
      8'b00111111: q[2] <= 9'b000101010;
      8'b01000000: q[2] <= 9'b000101010;
      8'b01000001: q[2] <= 9'b000101011;
      8'b01000010: q[2] <= 9'b000101100;
      8'b01000011: q[2] <= 9'b000101100;
      8'b01000100: q[2] <= 9'b000101101;
      8'b01000101: q[2] <= 9'b000101110;
      8'b01000110: q[2] <= 9'b000101110;
      8'b01000111: q[2] <= 9'b000101111;
      8'b01001000: q[2] <= 9'b000110000;
      8'b01001001: q[2] <= 9'b000110000;
      8'b01001010: q[2] <= 9'b000110001;
      8'b01001011: q[2] <= 9'b000110010;
      8'b01001100: q[2] <= 9'b000110010;
      8'b01001101: q[2] <= 9'b000110011;
      8'b01001110: q[2] <= 9'b000110100;
      8'b01001111: q[2] <= 9'b000110100;
      8'b01010000: q[2] <= 9'b000110101;
      8'b01010001: q[2] <= 9'b000110110;
      8'b01010010: q[2] <= 9'b000110110;
      8'b01010011: q[2] <= 9'b000110111;
      8'b01010100: q[2] <= 9'b000111000;
      8'b01010101: q[2] <= 9'b000111000;
      8'b01010110: q[2] <= 9'b000111001;
      8'b01010111: q[2] <= 9'b000111010;
      8'b01011000: q[2] <= 9'b000111010;
      8'b01011001: q[2] <= 9'b000111011;
      8'b01011010: q[2] <= 9'b000111100;
      8'b01011011: q[2] <= 9'b000111100;
      8'b01011100: q[2] <= 9'b000111101;
      8'b01011101: q[2] <= 9'b000111110;
      8'b01011110: q[2] <= 9'b000111110;
      8'b01011111: q[2] <= 9'b000111111;
      8'b01100000: q[2] <= 9'b001000000;
      8'b01100001: q[2] <= 9'b001000000;
      8'b01100010: q[2] <= 9'b001000001;
      8'b01100011: q[2] <= 9'b001000010;
      8'b01100100: q[2] <= 9'b001000010;
      8'b01100101: q[2] <= 9'b001000011;
      8'b01100110: q[2] <= 9'b001000100;
      8'b01100111: q[2] <= 9'b001000100;
      8'b01101000: q[2] <= 9'b001000101;
      8'b01101001: q[2] <= 9'b001000110;
      8'b01101010: q[2] <= 9'b001000110;
      8'b01101011: q[2] <= 9'b001000111;
      8'b01101100: q[2] <= 9'b001001000;
      8'b01101101: q[2] <= 9'b001001000;
      8'b01101110: q[2] <= 9'b001001001;
      8'b01101111: q[2] <= 9'b001001010;
      8'b01110000: q[2] <= 9'b001001010;
      8'b01110001: q[2] <= 9'b001001011;
      8'b01110010: q[2] <= 9'b001001100;
      8'b01110011: q[2] <= 9'b001001100;
      8'b01110100: q[2] <= 9'b001001101;
      8'b01110101: q[2] <= 9'b001001110;
      8'b01110110: q[2] <= 9'b001001110;
      8'b01110111: q[2] <= 9'b001001111;
      8'b01111000: q[2] <= 9'b001010000;
      8'b01111001: q[2] <= 9'b001010000;
      8'b01111010: q[2] <= 9'b001010001;
      8'b01111011: q[2] <= 9'b001010010;
      8'b01111100: q[2] <= 9'b001010010;
      8'b01111101: q[2] <= 9'b001010011;
      8'b01111110: q[2] <= 9'b001010100;
      8'b01111111: q[2] <= 9'b001010100;
      8'b10000000: q[2] <= 9'b001010101;
      8'b10000001: q[2] <= 9'b001010110;
      8'b10000010: q[2] <= 9'b001010110;
      8'b10000011: q[2] <= 9'b001010111;
      8'b10000100: q[2] <= 9'b001011000;
      8'b10000101: q[2] <= 9'b001011000;
      8'b10000110: q[2] <= 9'b001011001;
      8'b10000111: q[2] <= 9'b001011010;
      8'b10001000: q[2] <= 9'b001011010;
      8'b10001001: q[2] <= 9'b001011011;
      8'b10001010: q[2] <= 9'b001011100;
      8'b10001011: q[2] <= 9'b001011100;
      8'b10001100: q[2] <= 9'b001011101;
      8'b10001101: q[2] <= 9'b001011110;
      8'b10001110: q[2] <= 9'b001011110;
      8'b10001111: q[2] <= 9'b001011111;
      8'b10010000: q[2] <= 9'b001100000;
      8'b10010001: q[2] <= 9'b001100000;
      8'b10010010: q[2] <= 9'b001100001;
      8'b10010011: q[2] <= 9'b001100010;
      8'b10010100: q[2] <= 9'b001100010;
      8'b10010101: q[2] <= 9'b001100011;
      8'b10010110: q[2] <= 9'b001100100;
      8'b10010111: q[2] <= 9'b001100100;
      8'b10011000: q[2] <= 9'b001100101;
      8'b10011001: q[2] <= 9'b001100110;
      8'b10011010: q[2] <= 9'b001100110;
      8'b10011011: q[2] <= 9'b001100111;
      8'b10011100: q[2] <= 9'b001101000;
      8'b10011101: q[2] <= 9'b001101000;
      8'b10011110: q[2] <= 9'b001101001;
      8'b10011111: q[2] <= 9'b001101010;
      8'b10100000: q[2] <= 9'b001101010;
      8'b10100001: q[2] <= 9'b001101011;
      8'b10100010: q[2] <= 9'b001101100;
      8'b10100011: q[2] <= 9'b001101100;
      8'b10100100: q[2] <= 9'b001101101;
      8'b10100101: q[2] <= 9'b001101110;
      8'b10100110: q[2] <= 9'b001101110;
      8'b10100111: q[2] <= 9'b001101111;
      8'b10101000: q[2] <= 9'b001110000;
      8'b10101001: q[2] <= 9'b001110000;
      8'b10101010: q[2] <= 9'b001110001;
      8'b10101011: q[2] <= 9'b001110010;
      8'b10101100: q[2] <= 9'b001110010;
      8'b10101101: q[2] <= 9'b001110011;
      8'b10101110: q[2] <= 9'b001110100;
      8'b10101111: q[2] <= 9'b001110100;
      8'b10110000: q[2] <= 9'b001110101;
      8'b10110001: q[2] <= 9'b001110110;
      8'b10110010: q[2] <= 9'b001110110;
      8'b10110011: q[2] <= 9'b001110111;
      default: q[2] <= '0;
    endcase
    case (addr[7-1:0])
      7'b0000000: q[3] <= 9'b000000000;
      7'b0000001: q[3] <= 9'b000000000;
      7'b0000010: q[3] <= 9'b000000001;
      7'b0000011: q[3] <= 9'b000000001;
      7'b0000100: q[3] <= 9'b000000010;
      7'b0000101: q[3] <= 9'b000000010;
      7'b0000110: q[3] <= 9'b000000011;
      7'b0000111: q[3] <= 9'b000000011;
      7'b0001000: q[3] <= 9'b000000100;
      7'b0001001: q[3] <= 9'b000000100;
      7'b0001010: q[3] <= 9'b000000101;
      7'b0001011: q[3] <= 9'b000000101;
      7'b0001100: q[3] <= 9'b000000110;
      7'b0001101: q[3] <= 9'b000000110;
      7'b0001110: q[3] <= 9'b000000111;
      7'b0001111: q[3] <= 9'b000000111;
      7'b0010000: q[3] <= 9'b000001000;
      7'b0010001: q[3] <= 9'b000001000;
      7'b0010010: q[3] <= 9'b000001001;
      7'b0010011: q[3] <= 9'b000001001;
      7'b0010100: q[3] <= 9'b000001010;
      7'b0010101: q[3] <= 9'b000001010;
      7'b0010110: q[3] <= 9'b000001011;
      7'b0010111: q[3] <= 9'b000001011;
      7'b0011000: q[3] <= 9'b000001100;
      7'b0011001: q[3] <= 9'b000001100;
      7'b0011010: q[3] <= 9'b000001101;
      7'b0011011: q[3] <= 9'b000001101;
      7'b0011100: q[3] <= 9'b000001110;
      7'b0011101: q[3] <= 9'b000001110;
      7'b0011110: q[3] <= 9'b000001111;
      7'b0011111: q[3] <= 9'b000001111;
      7'b0100000: q[3] <= 9'b000010000;
      7'b0100001: q[3] <= 9'b000010000;
      7'b0100010: q[3] <= 9'b000010001;
      7'b0100011: q[3] <= 9'b000010001;
      7'b0100100: q[3] <= 9'b000010010;
      7'b0100101: q[3] <= 9'b000010010;
      7'b0100110: q[3] <= 9'b000010011;
      7'b0100111: q[3] <= 9'b000010011;
      7'b0101000: q[3] <= 9'b000010100;
      7'b0101001: q[3] <= 9'b000010100;
      7'b0101010: q[3] <= 9'b000010101;
      7'b0101011: q[3] <= 9'b000010101;
      7'b0101100: q[3] <= 9'b000010110;
      7'b0101101: q[3] <= 9'b000010110;
      7'b0101110: q[3] <= 9'b000010111;
      7'b0101111: q[3] <= 9'b000010111;
      7'b0110000: q[3] <= 9'b000011000;
      7'b0110001: q[3] <= 9'b000011000;
      7'b0110010: q[3] <= 9'b000011001;
      7'b0110011: q[3] <= 9'b000011001;
      7'b0110100: q[3] <= 9'b000011010;
      7'b0110101: q[3] <= 9'b000011010;
      7'b0110110: q[3] <= 9'b000011011;
      7'b0110111: q[3] <= 9'b000011011;
      7'b0111000: q[3] <= 9'b000011100;
      7'b0111001: q[3] <= 9'b000011100;
      7'b0111010: q[3] <= 9'b000011101;
      7'b0111011: q[3] <= 9'b000011101;
      7'b0111100: q[3] <= 9'b000011110;
      7'b0111101: q[3] <= 9'b000011110;
      7'b0111110: q[3] <= 9'b000011111;
      7'b0111111: q[3] <= 9'b000011111;
      7'b1000000: q[3] <= 9'b000100000;
      7'b1000001: q[3] <= 9'b000100000;
      7'b1000010: q[3] <= 9'b000100001;
      7'b1000011: q[3] <= 9'b000100001;
      7'b1000100: q[3] <= 9'b000100010;
      7'b1000101: q[3] <= 9'b000100010;
      7'b1000110: q[3] <= 9'b000100011;
      7'b1000111: q[3] <= 9'b000100011;
      7'b1001000: q[3] <= 9'b000100100;
      7'b1001001: q[3] <= 9'b000100100;
      7'b1001010: q[3] <= 9'b000100101;
      7'b1001011: q[3] <= 9'b000100101;
      7'b1001100: q[3] <= 9'b000100110;
      7'b1001101: q[3] <= 9'b000100110;
      7'b1001110: q[3] <= 9'b000100111;
      7'b1001111: q[3] <= 9'b000100111;
      7'b1010000: q[3] <= 9'b000101000;
      7'b1010001: q[3] <= 9'b000101000;
      7'b1010010: q[3] <= 9'b000101001;
      7'b1010011: q[3] <= 9'b000101001;
      7'b1010100: q[3] <= 9'b000101010;
      7'b1010101: q[3] <= 9'b000101010;
      7'b1010110: q[3] <= 9'b000101011;
      7'b1010111: q[3] <= 9'b000101011;
      7'b1011000: q[3] <= 9'b000101100;
      7'b1011001: q[3] <= 9'b000101100;
      7'b1011010: q[3] <= 9'b000101101;
      7'b1011011: q[3] <= 9'b000101101;
      7'b1011100: q[3] <= 9'b000101110;
      7'b1011101: q[3] <= 9'b000101110;
      7'b1011110: q[3] <= 9'b000101111;
      7'b1011111: q[3] <= 9'b000101111;
      7'b1100000: q[3] <= 9'b000110000;
      7'b1100001: q[3] <= 9'b000110000;
      7'b1100010: q[3] <= 9'b000110001;
      7'b1100011: q[3] <= 9'b000110001;
      7'b1100100: q[3] <= 9'b000110010;
      7'b1100101: q[3] <= 9'b000110010;
      7'b1100110: q[3] <= 9'b000110011;
      7'b1100111: q[3] <= 9'b000110011;
      7'b1101000: q[3] <= 9'b000110100;
      7'b1101001: q[3] <= 9'b000110100;
      7'b1101010: q[3] <= 9'b000110101;
      7'b1101011: q[3] <= 9'b000110101;
      7'b1101100: q[3] <= 9'b000110110;
      7'b1101101: q[3] <= 9'b000110110;
      7'b1101110: q[3] <= 9'b000110111;
      7'b1101111: q[3] <= 9'b000110111;
      7'b1110000: q[3] <= 9'b000111000;
      7'b1110001: q[3] <= 9'b000111000;
      7'b1110010: q[3] <= 9'b000111001;
      7'b1110011: q[3] <= 9'b000111001;
      7'b1110100: q[3] <= 9'b000111010;
      7'b1110101: q[3] <= 9'b000111010;
      7'b1110110: q[3] <= 9'b000111011;
      7'b1110111: q[3] <= 9'b000111011;
      default: q[3] <= '0;
    endcase
    case (addr[6-1:0])
      6'b000000: q[4] <= 9'b000000000;
      6'b000001: q[4] <= 9'b000000000;
      6'b000010: q[4] <= 9'b000000000;
      6'b000011: q[4] <= 9'b000000001;
      6'b000100: q[4] <= 9'b000000001;
      6'b000101: q[4] <= 9'b000000001;
      6'b000110: q[4] <= 9'b000000010;
      6'b000111: q[4] <= 9'b000000010;
      6'b001000: q[4] <= 9'b000000010;
      6'b001001: q[4] <= 9'b000000011;
      6'b001010: q[4] <= 9'b000000011;
      6'b001011: q[4] <= 9'b000000011;
      6'b001100: q[4] <= 9'b000000100;
      6'b001101: q[4] <= 9'b000000100;
      6'b001110: q[4] <= 9'b000000100;
      6'b001111: q[4] <= 9'b000000101;
      6'b010000: q[4] <= 9'b000000101;
      6'b010001: q[4] <= 9'b000000101;
      6'b010010: q[4] <= 9'b000000110;
      6'b010011: q[4] <= 9'b000000110;
      6'b010100: q[4] <= 9'b000000110;
      6'b010101: q[4] <= 9'b000000111;
      6'b010110: q[4] <= 9'b000000111;
      6'b010111: q[4] <= 9'b000000111;
      6'b011000: q[4] <= 9'b000001000;
      6'b011001: q[4] <= 9'b000001000;
      6'b011010: q[4] <= 9'b000001000;
      6'b011011: q[4] <= 9'b000001001;
      6'b011100: q[4] <= 9'b000001001;
      6'b011101: q[4] <= 9'b000001001;
      6'b011110: q[4] <= 9'b000001010;
      6'b011111: q[4] <= 9'b000001010;
      6'b100000: q[4] <= 9'b000001010;
      6'b100001: q[4] <= 9'b000001011;
      6'b100010: q[4] <= 9'b000001011;
      6'b100011: q[4] <= 9'b000001011;
      6'b100100: q[4] <= 9'b000001100;
      6'b100101: q[4] <= 9'b000001100;
      6'b100110: q[4] <= 9'b000001100;
      6'b100111: q[4] <= 9'b000001101;
      6'b101000: q[4] <= 9'b000001101;
      6'b101001: q[4] <= 9'b000001101;
      6'b101010: q[4] <= 9'b000001110;
      6'b101011: q[4] <= 9'b000001110;
      6'b101100: q[4] <= 9'b000001110;
      6'b101101: q[4] <= 9'b000001111;
      6'b101110: q[4] <= 9'b000001111;
      6'b101111: q[4] <= 9'b000001111;
      6'b110000: q[4] <= 9'b000010000;
      6'b110001: q[4] <= 9'b000010000;
      6'b110010: q[4] <= 9'b000010000;
      6'b110011: q[4] <= 9'b000010001;
      6'b110100: q[4] <= 9'b000010001;
      6'b110101: q[4] <= 9'b000010001;
      6'b110110: q[4] <= 9'b000010010;
      6'b110111: q[4] <= 9'b000010010;
      6'b111000: q[4] <= 9'b000010010;
      6'b111001: q[4] <= 9'b000010011;
      6'b111010: q[4] <= 9'b000010011;
      6'b111011: q[4] <= 9'b000010011;
      default: q[4] <= '0;
    endcase
  end

  assign addrOut = scaleNum<5?q[scaleNum]:'1
endmodule
