module heu_sum_lut
  (
    /*
     * Inputs
     */
    input [8:0] d,

    /*
     * Outputs
     */
    output reg [7:0] q
  );

  always_comb begin
    case (d)
      9'b000000000: q <= 8'b00000000;
      9'b000000001: q <= 8'b00000000;
      9'b000000010: q <= 8'b00000001;
      9'b000000011: q <= 8'b00000001;
      9'b000000100: q <= 8'b00000010;
      9'b000000101: q <= 8'b00000011;
      9'b000000110: q <= 8'b00000011;
      9'b000000111: q <= 8'b00000100;
      9'b000001000: q <= 8'b00000101;
      9'b000001001: q <= 8'b00000101;
      9'b000001010: q <= 8'b00000110;
      9'b000001011: q <= 8'b00000111;
      9'b000001100: q <= 8'b00000111;
      9'b000001101: q <= 8'b00001000;
      9'b000001110: q <= 8'b00001000;
      9'b000001111: q <= 8'b00001001;
      9'b000010000: q <= 8'b00001010;
      9'b000010001: q <= 8'b00001010;
      9'b000010010: q <= 8'b00001011;
      9'b000010011: q <= 8'b00001100;
      9'b000010100: q <= 8'b00001100;
      9'b000010101: q <= 8'b00001101;
      9'b000010110: q <= 8'b00001110;
      9'b000010111: q <= 8'b00001110;
      9'b000011000: q <= 8'b00001111;
      9'b000011001: q <= 8'b00001111;
      9'b000011010: q <= 8'b00010000;
      9'b000011011: q <= 8'b00010001;
      9'b000011100: q <= 8'b00010001;
      9'b000011101: q <= 8'b00010010;
      9'b000011110: q <= 8'b00010011;
      9'b000011111: q <= 8'b00010011;
      9'b000100000: q <= 8'b00010100;
      9'b000100001: q <= 8'b00010101;
      9'b000100010: q <= 8'b00010101;
      9'b000100011: q <= 8'b00010110;
      9'b000100100: q <= 8'b00010110;
      9'b000100101: q <= 8'b00010111;
      9'b000100110: q <= 8'b00011000;
      9'b000100111: q <= 8'b00011000;
      9'b000101000: q <= 8'b00011001;
      9'b000101001: q <= 8'b00011010;
      9'b000101010: q <= 8'b00011010;
      9'b000101011: q <= 8'b00011011;
      9'b000101100: q <= 8'b00011100;
      9'b000101101: q <= 8'b00011100;
      9'b000101110: q <= 8'b00011101;
      9'b000101111: q <= 8'b00011101;
      9'b000110000: q <= 8'b00011110;
      9'b000110001: q <= 8'b00011111;
      9'b000110010: q <= 8'b00011111;
      9'b000110011: q <= 8'b00100000;
      9'b000110100: q <= 8'b00100001;
      9'b000110101: q <= 8'b00100001;
      9'b000110110: q <= 8'b00100010;
      9'b000110111: q <= 8'b00100011;
      9'b000111000: q <= 8'b00100011;
      9'b000111001: q <= 8'b00100100;
      9'b000111010: q <= 8'b00100100;
      9'b000111011: q <= 8'b00100101;
      9'b000111100: q <= 8'b00100110;
      9'b000111101: q <= 8'b00100110;
      9'b000111110: q <= 8'b00100111;
      9'b000111111: q <= 8'b00101000;
      9'b001000000: q <= 8'b00101000;
      9'b001000001: q <= 8'b00101001;
      9'b001000010: q <= 8'b00101010;
      9'b001000011: q <= 8'b00101010;
      9'b001000100: q <= 8'b00101011;
      9'b001000101: q <= 8'b00101011;
      9'b001000110: q <= 8'b00101100;
      9'b001000111: q <= 8'b00101101;
      9'b001001000: q <= 8'b00101101;
      9'b001001001: q <= 8'b00101110;
      9'b001001010: q <= 8'b00101111;
      9'b001001011: q <= 8'b00101111;
      9'b001001100: q <= 8'b00110000;
      9'b001001101: q <= 8'b00110001;
      9'b001001110: q <= 8'b00110001;
      9'b001001111: q <= 8'b00110010;
      9'b001010000: q <= 8'b00110011;
      9'b001010001: q <= 8'b00110011;
      9'b001010010: q <= 8'b00110100;
      9'b001010011: q <= 8'b00110100;
      9'b001010100: q <= 8'b00110101;
      9'b001010101: q <= 8'b00110110;
      9'b001010110: q <= 8'b00110110;
      9'b001010111: q <= 8'b00110111;
      9'b001011000: q <= 8'b00111000;
      9'b001011001: q <= 8'b00111000;
      9'b001011010: q <= 8'b00111001;
      9'b001011011: q <= 8'b00111010;
      9'b001011100: q <= 8'b00111010;
      9'b001011101: q <= 8'b00111011;
      9'b001011110: q <= 8'b00111011;
      9'b001011111: q <= 8'b00111100;
      9'b001100000: q <= 8'b00111101;
      9'b001100001: q <= 8'b00111101;
      9'b001100010: q <= 8'b00111110;
      9'b001100011: q <= 8'b00111111;
      9'b001100100: q <= 8'b00111111;
      9'b001100101: q <= 8'b01000000;
      9'b001100110: q <= 8'b01000001;
      9'b001100111: q <= 8'b01000001;
      9'b001101000: q <= 8'b01000010;
      9'b001101001: q <= 8'b01000010;
      9'b001101010: q <= 8'b01000011;
      9'b001101011: q <= 8'b01000100;
      9'b001101100: q <= 8'b01000100;
      9'b001101101: q <= 8'b01000101;
      9'b001101110: q <= 8'b01000110;
      9'b001101111: q <= 8'b01000110;
      9'b001110000: q <= 8'b01000111;
      9'b001110001: q <= 8'b01001000;
      9'b001110010: q <= 8'b01001000;
      9'b001110011: q <= 8'b01001001;
      9'b001110100: q <= 8'b01001001;
      9'b001110101: q <= 8'b01001010;
      9'b001110110: q <= 8'b01001011;
      9'b001110111: q <= 8'b01001011;
      9'b001111000: q <= 8'b01001100;
      9'b001111001: q <= 8'b01001101;
      9'b001111010: q <= 8'b01001101;
      9'b001111011: q <= 8'b01001110;
      9'b001111100: q <= 8'b01001111;
      9'b001111101: q <= 8'b01001111;
      9'b001111110: q <= 8'b01010000;
      9'b001111111: q <= 8'b01010000;
      9'b010000000: q <= 8'b01010001;
      9'b010000001: q <= 8'b01010010;
      9'b010000010: q <= 8'b01010010;
      9'b010000011: q <= 8'b01010011;
      9'b010000100: q <= 8'b01010100;
      9'b010000101: q <= 8'b01010100;
      9'b010000110: q <= 8'b01010101;
      9'b010000111: q <= 8'b01010110;
      9'b010001000: q <= 8'b01010110;
      9'b010001001: q <= 8'b01010111;
      9'b010001010: q <= 8'b01010111;
      9'b010001011: q <= 8'b01011000;
      9'b010001100: q <= 8'b01011001;
      9'b010001101: q <= 8'b01011001;
      9'b010001110: q <= 8'b01011010;
      9'b010001111: q <= 8'b01011011;
      9'b010010000: q <= 8'b01011011;
      9'b010010001: q <= 8'b01011100;
      9'b010010010: q <= 8'b01011101;
      9'b010010011: q <= 8'b01011101;
      9'b010010100: q <= 8'b01011110;
      9'b010010101: q <= 8'b01011110;
      9'b010010110: q <= 8'b01011111;
      9'b010010111: q <= 8'b01100000;
      9'b010011000: q <= 8'b01100000;
      9'b010011001: q <= 8'b01100001;
      9'b010011010: q <= 8'b01100010;
      9'b010011011: q <= 8'b01100010;
      9'b010011100: q <= 8'b01100011;
      9'b010011101: q <= 8'b01100100;
      9'b010011110: q <= 8'b01100100;
      9'b010011111: q <= 8'b01100101;
      9'b010100000: q <= 8'b01100110;
      9'b010100001: q <= 8'b01100110;
      9'b010100010: q <= 8'b01100111;
      9'b010100011: q <= 8'b01100111;
      9'b010100100: q <= 8'b01101000;
      9'b010100101: q <= 8'b01101001;
      9'b010100110: q <= 8'b01101001;
      9'b010100111: q <= 8'b01101010;
      9'b010101000: q <= 8'b01101011;
      9'b010101001: q <= 8'b01101011;
      9'b010101010: q <= 8'b01101100;
      9'b010101011: q <= 8'b01101101;
      9'b010101100: q <= 8'b01101101;
      9'b010101101: q <= 8'b01101110;
      9'b010101110: q <= 8'b01101110;
      9'b010101111: q <= 8'b01101111;
      9'b010110000: q <= 8'b01110000;
      9'b010110001: q <= 8'b01110000;
      9'b010110010: q <= 8'b01110001;
      9'b010110011: q <= 8'b01110010;
      9'b010110100: q <= 8'b01110010;
      9'b010110101: q <= 8'b01110011;
      9'b010110110: q <= 8'b01110100;
      9'b010110111: q <= 8'b01110100;
      9'b010111000: q <= 8'b01110101;
      9'b010111001: q <= 8'b01110101;
      9'b010111010: q <= 8'b01110110;
      9'b010111011: q <= 8'b01110111;
      9'b010111100: q <= 8'b01110111;
      9'b010111101: q <= 8'b01111000;
      9'b010111110: q <= 8'b01111001;
      9'b010111111: q <= 8'b01111001;
      9'b011000000: q <= 8'b01111010;
      9'b011000001: q <= 8'b01111011;
      9'b011000010: q <= 8'b01111011;
      9'b011000011: q <= 8'b01111100;
      9'b011000100: q <= 8'b01111100;
      9'b011000101: q <= 8'b01111101;
      9'b011000110: q <= 8'b01111110;
      9'b011000111: q <= 8'b01111110;
      9'b011001000: q <= 8'b01111111;
      9'b011001001: q <= 8'b10000000;
      9'b011001010: q <= 8'b10000000;
      9'b011001011: q <= 8'b10000001;
      9'b011001100: q <= 8'b10000010;
      9'b011001101: q <= 8'b10000010;
      9'b011001110: q <= 8'b10000011;
      9'b011001111: q <= 8'b10000011;
      9'b011010000: q <= 8'b10000100;
      9'b011010001: q <= 8'b10000101;
      9'b011010010: q <= 8'b10000101;
      9'b011010011: q <= 8'b10000110;
      9'b011010100: q <= 8'b10000111;
      9'b011010101: q <= 8'b10000111;
      9'b011010110: q <= 8'b10001000;
      9'b011010111: q <= 8'b10001001;
      9'b011011000: q <= 8'b10001001;
      9'b011011001: q <= 8'b10001010;
      9'b011011010: q <= 8'b10001010;
      9'b011011011: q <= 8'b10001011;
      9'b011011100: q <= 8'b10001100;
      9'b011011101: q <= 8'b10001100;
      9'b011011110: q <= 8'b10001101;
      9'b011011111: q <= 8'b10001110;
      9'b011100000: q <= 8'b10001110;
      9'b011100001: q <= 8'b10001111;
      9'b011100010: q <= 8'b10010000;
      9'b011100011: q <= 8'b10010000;
      9'b011100100: q <= 8'b10010001;
      9'b011100101: q <= 8'b10010001;
      9'b011100110: q <= 8'b10010010;
      9'b011100111: q <= 8'b10010011;
      9'b011101000: q <= 8'b10010011;
      9'b011101001: q <= 8'b10010100;
      9'b011101010: q <= 8'b10010101;
      9'b011101011: q <= 8'b10010101;
      9'b011101100: q <= 8'b10010110;
      9'b011101101: q <= 8'b10010111;
      9'b011101110: q <= 8'b10010111;
      9'b011101111: q <= 8'b10011000;
      9'b011110000: q <= 8'b10011001;
      9'b011110001: q <= 8'b10011001;
      9'b011110010: q <= 8'b10011010;
      9'b011110011: q <= 8'b10011010;
      9'b011110100: q <= 8'b10011011;
      9'b011110101: q <= 8'b10011100;
      9'b011110110: q <= 8'b10011100;
      9'b011110111: q <= 8'b10011101;
      9'b011111000: q <= 8'b10011110;
      9'b011111001: q <= 8'b10011110;
      9'b011111010: q <= 8'b10011111;
      9'b011111011: q <= 8'b10100000;
      9'b011111100: q <= 8'b10100000;
      9'b011111101: q <= 8'b10100001;
      9'b011111110: q <= 8'b10100001;
      9'b011111111: q <= 8'b10100010;
      9'b100000000: q <= 8'b10100011;
      9'b100000001: q <= 8'b10100011;
      9'b100000010: q <= 8'b10100100;
      9'b100000011: q <= 8'b10100101;
      9'b100000100: q <= 8'b10100101;
      9'b100000101: q <= 8'b10100110;
      9'b100000110: q <= 8'b10100111;
      9'b100000111: q <= 8'b10100111;
      9'b100001000: q <= 8'b10101000;
      9'b100001001: q <= 8'b10101000;
      9'b100001010: q <= 8'b10101001;
      9'b100001011: q <= 8'b10101010;
      9'b100001100: q <= 8'b10101010;
      9'b100001101: q <= 8'b10101011;
      9'b100001110: q <= 8'b10101100;
      9'b100001111: q <= 8'b10101100;
      9'b100010000: q <= 8'b10101101;
      9'b100010001: q <= 8'b10101110;
      9'b100010010: q <= 8'b10101110;
      9'b100010011: q <= 8'b10101111;
      9'b100010100: q <= 8'b10101111;
      9'b100010101: q <= 8'b10110000;
      9'b100010110: q <= 8'b10110001;
      9'b100010111: q <= 8'b10110001;
      9'b100011000: q <= 8'b10110010;
      9'b100011001: q <= 8'b10110011;
      9'b100011010: q <= 8'b10110011;
      9'b100011011: q <= 8'b10110100;
      9'b100011100: q <= 8'b10110101;
      9'b100011101: q <= 8'b10110101;
      9'b100011110: q <= 8'b10110110;
      9'b100011111: q <= 8'b10110110;
      9'b100100000: q <= 8'b10110111;
      9'b100100001: q <= 8'b10111000;
      9'b100100010: q <= 8'b10111000;
      9'b100100011: q <= 8'b10111001;
      9'b100100100: q <= 8'b10111010;
      9'b100100101: q <= 8'b10111010;
      9'b100100110: q <= 8'b10111011;
      9'b100100111: q <= 8'b10111100;
      9'b100101000: q <= 8'b10111100;
      9'b100101001: q <= 8'b10111101;
      9'b100101010: q <= 8'b10111101;
      9'b100101011: q <= 8'b10111110;
      9'b100101100: q <= 8'b10111111;
      9'b100101101: q <= 8'b10111111;
      9'b100101110: q <= 8'b11000000;
      9'b100101111: q <= 8'b11000001;
      9'b100110000: q <= 8'b11000001;
      9'b100110001: q <= 8'b11000010;
      9'b100110010: q <= 8'b11000011;
      9'b100110011: q <= 8'b11000011;
      9'b100110100: q <= 8'b11000100;
      9'b100110101: q <= 8'b11000100;
      9'b100110110: q <= 8'b11000101;
      9'b100110111: q <= 8'b11000110;
      9'b100111000: q <= 8'b11000110;
      9'b100111001: q <= 8'b11000111;
      9'b100111010: q <= 8'b11001000;
      9'b100111011: q <= 8'b11001000;
      9'b100111100: q <= 8'b11001001;
      9'b100111101: q <= 8'b11001010;
      9'b100111110: q <= 8'b11001010;
      9'b100111111: q <= 8'b11001011;
      9'b101000000: q <= 8'b11001100;
      9'b101000001: q <= 8'b11001100;
      9'b101000010: q <= 8'b11001101;
      9'b101000011: q <= 8'b11001101;
      9'b101000100: q <= 8'b11001110;
      9'b101000101: q <= 8'b11001111;
      9'b101000110: q <= 8'b11001111;
      9'b101000111: q <= 8'b11010000;
      9'b101001000: q <= 8'b11010001;
      9'b101001001: q <= 8'b11010001;
      9'b101001010: q <= 8'b11010010;
      9'b101001011: q <= 8'b11010011;
      9'b101001100: q <= 8'b11010011;
      9'b101001101: q <= 8'b11010100;
      9'b101001110: q <= 8'b11010100;
      9'b101001111: q <= 8'b11010101;
      9'b101010000: q <= 8'b11010110;
      9'b101010001: q <= 8'b11010110;
      9'b101010010: q <= 8'b11010111;
      9'b101010011: q <= 8'b11011000;
      9'b101010100: q <= 8'b11011000;
      9'b101010101: q <= 8'b11011001;
      9'b101010110: q <= 8'b11011010;
      9'b101010111: q <= 8'b11011010;
      9'b101011000: q <= 8'b11011011;
      9'b101011001: q <= 8'b11011011;
      9'b101011010: q <= 8'b11011100;
      9'b101011011: q <= 8'b11011101;
      9'b101011100: q <= 8'b11011101;
      9'b101011101: q <= 8'b11011110;
      9'b101011110: q <= 8'b11011111;
      9'b101011111: q <= 8'b11011111;
      9'b101100000: q <= 8'b11100000;
      9'b101100001: q <= 8'b11100001;
      9'b101100010: q <= 8'b11100001;
      9'b101100011: q <= 8'b11100010;
      9'b101100100: q <= 8'b11100010;
      9'b101100101: q <= 8'b11100011;
      9'b101100110: q <= 8'b11100100;
      9'b101100111: q <= 8'b11100100;
      9'b101101000: q <= 8'b11100101;
      9'b101101001: q <= 8'b11100110;
      9'b101101010: q <= 8'b11100110;
      9'b101101011: q <= 8'b11100111;
      9'b101101100: q <= 8'b11101000;
      9'b101101101: q <= 8'b11101000;
      9'b101101110: q <= 8'b11101001;
      9'b101101111: q <= 8'b11101001;
      9'b101110000: q <= 8'b11101010;
      9'b101110001: q <= 8'b11101011;
      9'b101110010: q <= 8'b11101011;
      9'b101110011: q <= 8'b11101100;
      9'b101110100: q <= 8'b11101101;
      9'b101110101: q <= 8'b11101101;
      9'b101110110: q <= 8'b11101110;
      9'b101110111: q <= 8'b11101111;
      9'b101111000: q <= 8'b11101111;
      9'b101111001: q <= 8'b11110000;
      9'b101111010: q <= 8'b11110000;
      9'b101111011: q <= 8'b11110001;
      9'b101111100: q <= 8'b11110010;
      9'b101111101: q <= 8'b11110010;
      9'b101111110: q <= 8'b11110011;
      9'b101111111: q <= 8'b11110100;
      9'b110000000: q <= 8'b11110100;
      9'b110000001: q <= 8'b11110101;
      9'b110000010: q <= 8'b11110110;
      9'b110000011: q <= 8'b11110110;
      9'b110000100: q <= 8'b11110111;
      9'b110000101: q <= 8'b11110111;
      9'b110000110: q <= 8'b11111000;
      9'b110000111: q <= 8'b11111001;
      9'b110001000: q <= 8'b11111001;
      9'b110001001: q <= 8'b11111010;
      9'b110001010: q <= 8'b11111011;
      9'b110001011: q <= 8'b11111011;
      9'b110001100: q <= 8'b11111100;
      9'b110001101: q <= 8'b11111101;
      9'b110001110: q <= 8'b11111101;
      9'b110001111: q <= 8'b11111110;
      9'b110010000: q <= 8'b11111111;
      default: q <= 0;
    endcase
  end

endmodule
