

module ccip_mmio (
    input pClk,
    
  );
